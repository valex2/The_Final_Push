module wave_display_tb (

);

endmodule