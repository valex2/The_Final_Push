module wave_capture_tb (

);

endmodule